// 이곳에 1차과제 제출물이 들어갈 전체 Main 모듈 작성