module SNN(
    input logic clk,
    input logic reset
);


endmodule